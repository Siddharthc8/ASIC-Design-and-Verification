class async_fifo_common extends uvm_component;


endclass