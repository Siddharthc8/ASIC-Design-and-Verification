
// typedef uvm_sequencer#(write_tx) write_sqr;

class write_sqr extends uvm_sequencer#(write_tx);
`uvm_component_utils(write_sqr)

    `NEW_COMP

endclass