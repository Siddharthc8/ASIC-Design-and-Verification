// typedef uvm_sequencer#(read_tx) read_sqr;

class read_sqr extends uvm_sequencer#(read_tx);
`uvm_component_utils(read_sqr)

    `NEW_COMP

endclass