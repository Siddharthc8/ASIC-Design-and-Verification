interface axi_intf(input bit aclk, arst);


endinterface